module fsm(Strobe, RW, M, V, CtrSig, LdCtr, RdyEn, Rdy, W, MStrobe, MRW, Wsel, RSel);
	
	input logic Strobe;
	input logic RW
	input logic M
	input logic V
	input logic CtrSig
	
	output logic LdCtr
	output logic RdyEn
	output logic Rdy
	output logic W 
	output logic MStrobe
	output logic MRW
	output logic RSel
	
	parameter [3:0] S0 = 4'd0,
     S1 = 4'd1,
     S2 = 4'd2,
     S3 = 4'd3,
     S4 = 4'd4,
     S5 = 4'd5,
     S6 = 4'd6,
     S7 = 4'd7,
	 s8 = 4'd8,
	 s9 = 4'd9,
     Idle = 4'd10;

   logic [3:0] CURRENT_STATE;
   logic [3:0] NEXT_STATE;
   //past this point is merely copy/pasted 
   

   always @(CURRENT_STATE or Strobe)
     begin
 	case(CURRENT_STATE)
	  Idle:	
	    if (Strobe == 1'b0)
	      begin
		 LdCtr = 1'b1;
		 RdyEn = 1'b0;
		 Rdy   = 1'b0;
		 NEXT_STATE <=  Idle;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S0;
	      end
	  
	  S0:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b0;
		 NEXT_STATE <=  S1;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S0;
	      end	
	  
	  S1:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b0;
		 NEXT_STATE <=  Idle;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S2;
	      end	

	  S2:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b0;
		 NEXT_STATE <=  S1;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S3;
	      end	

	  S3:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b0;
		 NEXT_STATE <=  S4;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S0;
	      end	

	  S4:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b0;
		 NEXT_STATE <=  Idle;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S5;
	      end	

	  S5:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b0;
		 NEXT_STATE <=  S1;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S6;
	      end	

	  S6:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b0;
		 NEXT_STATE <=  S7;
	      end else begin
		 Z = 1'b0;
		 NEXT_STATE <=  S0;
	      end	

	  S7:	
	    if (X == 1'b0)
	      begin
		 Z = 1'b1;
		 NEXT_STATE <=  Idle;
	      end else begin
		 Z = 1'b1;
		 NEXT_STATE <=  S5;
	      end
	  
	  s8:
		if
		  end
	  s9:
		  end
	  
	  default: 
	    begin
	       NEXT_STATE <=  S0;
	       Z = 1'b0;	     
	    end
	  
	endcase // case (CURRENT_STATE)	
     end // always @ (CURRENT_STATE or X)

endmodule //fsm